// Code your design here
`include "sram.v"
`include "apb_slave.v"